module top;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import pkg_lib::*;
    initial run_test("txn_test");
endmodule
