package pkg_lib;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    typedef class txn;

    // Typdefs
    typedef txn q_of_txn_t[$];
    typedef int q_of_idx[$];

    // Items
    `include "txn.sv"

    // Agent
    typedef uvm_sequencer #(txn) txn_sqr;
    `include "txn_drv.sv"
    `include "seq_lib.sv"

    // Callbacks
   `include "txn_callbacks.sv"

    // Components
    `include "txn_route.sv"
    `include "ooo_comparator.sv"
    `include "txn_ooo_comp.sv"

    // Tests
    `include "test_lib.sv"

endpackage
